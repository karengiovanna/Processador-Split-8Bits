library ieee;
use ieee.std_logic_1164.all;

entity multiplexador_banco_ula is 
    port(
        ula_src : in std_logic;
        dado_lido  
    );
end multiplexador_banco_ula;

architecture multiplexador_comportamento of multiplexador_banco_ula
    begin
        
    end multiplexador_comportamento;
